//top level module for single cycle CPU
//makes all interconnections between different
//processing blocks

module CPU_single();

	
	//instantiate all wires here
	
	
	
	//program counter goes here
	//PC module
	
	//CPU control unit
	
	//ALU control unit
	
	//regfile instantiation
	
	//ALU instantiation
	
	//LSR, LSL instruction support here
	
	
	




endmodule 